-------------------------------------------------------------------------------
-- Title      : negative disparity rom
-- Project    : 
-------------------------------------------------------------------------------
-- File       : enc_8_10_rom2p.vhd
-- Author     : amr  <amr@laptop>
-- Company    : 
-- Created    : 2014-10-15
-- Last update: 24-10-2014
-- Platform   : 
-- Standard   : VHDL'87
-------------------------------------------------------------------------------
-- Description: a negative disparity rom
-------------------------------------------------------------------------------
-- Copyright (c) 2014 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2014-10-15  1.0      amr     Created
-------------------------------------------------------------------------------
library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

entity enc_8_10_rom2p is
  
  port (
    clk       : in  std_logic;
    address_a : in  std_logic_vector(8 downto 0);
    address_b : in  std_logic_vector(8 downto 0);
    rde_a     : in  std_logic;
    rde_b     : in  std_logic;
    dout_a    : out std_logic_vector(19 downto 0);
    dout_b    : out std_logic_vector(19 downto 0)
    );


end enc_8_10_rom2p;


architecture behav of enc_8_10_rom2p is

  type ROM_t is array (0 to 267) of std_logic_vector(19 downto 0);
  shared variable aRAM : ROM_t := (

    "10" & x"74" & "01" & x"8b",
    "01" & x"d4" & "10" & x"2b",
    "10" & x"d4" & "01" & x"2b",
    "11" & x"1b" & "11" & x"14",
    "11" & x"54" & "00" & x"ab",
    "10" & x"9b" & "10" & x"94",
    "01" & x"9b" & "01" & x"94",
    "11" & x"8b" & "00" & x"74",
    "11" & x"94" & "00" & x"6b",
    "10" & x"5b" & "10" & x"54",
    "01" & x"5b" & "01" & x"54",
    "11" & x"4b" & "11" & x"44",
    "00" & x"db" & "00" & x"d4",
    "10" & x"cb" & "10" & x"c4",
    "01" & x"cb" & "01" & x"c4",
    "01" & x"74" & "10" & x"8b",
    "01" & x"b4" & "10" & x"4b",
    "10" & x"3b" & "10" & x"34",
    "01" & x"3b" & "01" & x"34",
    "11" & x"2b" & "11" & x"24",
    "00" & x"bb" & "00" & x"b4",
    "10" & x"ab" & "10" & x"a4",
    "01" & x"ab" & "01" & x"a4",
    "11" & x"a4" & "00" & x"5b",
    "11" & x"34" & "00" & x"cb",
    "10" & x"6b" & "10" & x"64",
    "01" & x"6b" & "01" & x"64",
    "11" & x"64" & "00" & x"9b",
    "00" & x"eb" & "00" & x"e4",
    "10" & x"e4" & "01" & x"1b",
    "01" & x"e4" & "10" & x"1b",
    "10" & x"b4" & "01" & x"4b",
    "10" & x"79" & "01" & x"89",
    "01" & x"d9" & "10" & x"29",
    "10" & x"d9" & "01" & x"29",
    "11" & x"19" & "11" & x"19",
    "11" & x"59" & "00" & x"a9",
    "10" & x"99" & "10" & x"99",
    "01" & x"99" & "01" & x"99",
    "11" & x"89" & "00" & x"79",
    "11" & x"99" & "00" & x"69",
    "10" & x"59" & "10" & x"59",
    "01" & x"59" & "01" & x"59",
    "11" & x"49" & "11" & x"49",
    "00" & x"d9" & "00" & x"d9",
    "10" & x"c9" & "10" & x"c9",
    "01" & x"c9" & "01" & x"c9",
    "01" & x"79" & "10" & x"89",
    "01" & x"b9" & "10" & x"49",
    "10" & x"39" & "10" & x"39",
    "01" & x"39" & "01" & x"39",
    "11" & x"29" & "11" & x"29",
    "00" & x"b9" & "00" & x"b9",
    "10" & x"a9" & "10" & x"a9",
    "01" & x"a9" & "01" & x"a9",
    "11" & x"a9" & "00" & x"59",
    "11" & x"39" & "00" & x"c9",
    "10" & x"69" & "10" & x"69",
    "01" & x"69" & "01" & x"69",
    "11" & x"69" & "00" & x"99",
    "00" & x"e9" & "00" & x"e9",
    "10" & x"e9" & "01" & x"19",
    "01" & x"e9" & "10" & x"19",
    "10" & x"b9" & "01" & x"49",
    "10" & x"75" & "01" & x"85",
    "01" & x"d5" & "10" & x"25",
    "10" & x"d5" & "01" & x"25",
    "11" & x"15" & "11" & x"15",
    "11" & x"55" & "00" & x"a5",
    "10" & x"95" & "10" & x"95",
    "01" & x"95" & "01" & x"95",
    "11" & x"85" & "00" & x"75",
    "11" & x"95" & "00" & x"65",
    "10" & x"55" & "10" & x"55",
    "01" & x"55" & "01" & x"55",
    "11" & x"45" & "11" & x"45",
    "00" & x"d5" & "00" & x"d5",
    "10" & x"c5" & "10" & x"c5",
    "01" & x"c5" & "01" & x"c5",
    "01" & x"75" & "10" & x"85",
    "01" & x"b5" & "10" & x"45",
    "10" & x"35" & "10" & x"35",
    "01" & x"35" & "01" & x"35",
    "11" & x"25" & "11" & x"25",
    "00" & x"b5" & "00" & x"b5",
    "10" & x"a5" & "10" & x"a5",
    "01" & x"a5" & "01" & x"a5",
    "11" & x"a5" & "00" & x"55",
    "11" & x"35" & "00" & x"c5",
    "10" & x"65" & "10" & x"65",
    "01" & x"65" & "01" & x"65",
    "11" & x"65" & "00" & x"95",
    "00" & x"e5" & "00" & x"e5",
    "10" & x"e5" & "01" & x"15",
    "01" & x"e5" & "10" & x"15",
    "10" & x"b5" & "01" & x"45",
    "10" & x"73" & "01" & x"8c",
    "01" & x"d3" & "10" & x"2c",
    "10" & x"d3" & "01" & x"2c",
    "11" & x"1c" & "11" & x"13",
    "11" & x"53" & "00" & x"ac",
    "10" & x"9c" & "10" & x"93",
    "01" & x"9c" & "01" & x"93",
    "11" & x"8c" & "00" & x"73",
    "11" & x"93" & "00" & x"6c",
    "10" & x"5c" & "10" & x"53",
    "01" & x"5c" & "01" & x"53",
    "11" & x"4c" & "11" & x"43",
    "00" & x"dc" & "00" & x"d3",
    "10" & x"cc" & "10" & x"c3",
    "01" & x"cc" & "01" & x"c3",
    "01" & x"73" & "10" & x"8c",
    "01" & x"b3" & "10" & x"4c",
    "10" & x"3c" & "10" & x"33",
    "01" & x"3c" & "01" & x"33",
    "11" & x"2c" & "11" & x"23",
    "00" & x"bc" & "00" & x"b3",
    "10" & x"ac" & "10" & x"a3",
    "01" & x"ac" & "01" & x"a3",
    "11" & x"a3" & "00" & x"5c",
    "11" & x"33" & "00" & x"cc",
    "10" & x"6c" & "10" & x"63",
    "01" & x"6c" & "01" & x"63",
    "11" & x"63" & "00" & x"9c",
    "00" & x"ec" & "00" & x"e3",
    "10" & x"e3" & "01" & x"1c",
    "01" & x"e3" & "10" & x"1c",
    "10" & x"b3" & "01" & x"4c",
    "10" & x"72" & "01" & x"8d",
    "01" & x"d2" & "10" & x"2d",
    "10" & x"d2" & "01" & x"2d",
    "11" & x"1d" & "11" & x"12",
    "11" & x"52" & "00" & x"ad",
    "10" & x"9d" & "10" & x"92",
    "01" & x"9d" & "01" & x"92",
    "11" & x"8d" & "00" & x"72",
    "11" & x"92" & "00" & x"6d",
    "10" & x"5d" & "10" & x"52",
    "01" & x"5d" & "01" & x"52",
    "11" & x"4d" & "11" & x"42",
    "00" & x"dd" & "00" & x"d2",
    "10" & x"cd" & "10" & x"c2",
    "01" & x"cd" & "01" & x"c2",
    "01" & x"72" & "10" & x"8d",
    "01" & x"b2" & "10" & x"4d",
    "10" & x"3d" & "10" & x"32",
    "01" & x"3d" & "01" & x"32",
    "11" & x"2d" & "11" & x"22",
    "00" & x"bd" & "00" & x"b2",
    "10" & x"ad" & "10" & x"a2",
    "01" & x"ad" & "01" & x"a2",
    "11" & x"a2" & "00" & x"5d",
    "11" & x"32" & "00" & x"cd",
    "10" & x"6d" & "10" & x"62",
    "01" & x"6d" & "01" & x"62",
    "11" & x"62" & "00" & x"9d",
    "00" & x"ed" & "00" & x"e2",
    "10" & x"e2" & "01" & x"1d",
    "01" & x"e2" & "10" & x"1d",
    "10" & x"b2" & "01" & x"4d",
    "10" & x"7a" & "01" & x"8a",
    "01" & x"da" & "10" & x"2a",
    "10" & x"da" & "01" & x"2a",
    "11" & x"1a" & "11" & x"1a",
    "11" & x"5a" & "00" & x"aa",
    "10" & x"9a" & "10" & x"9a",
    "01" & x"9a" & "01" & x"9a",
    "11" & x"8a" & "00" & x"7a",
    "11" & x"9a" & "00" & x"6a",
    "10" & x"5a" & "10" & x"5a",
    "01" & x"5a" & "01" & x"5a",
    "11" & x"4a" & "11" & x"4a",
    "00" & x"da" & "00" & x"da",
    "10" & x"ca" & "10" & x"ca",
    "01" & x"ca" & "01" & x"ca",
    "01" & x"7a" & "10" & x"8a",
    "01" & x"ba" & "10" & x"4a",
    "10" & x"3a" & "10" & x"3a",
    "01" & x"3a" & "01" & x"3a",
    "11" & x"2a" & "11" & x"2a",
    "00" & x"ba" & "00" & x"ba",
    "10" & x"aa" & "10" & x"aa",
    "01" & x"aa" & "01" & x"aa",
    "11" & x"aa" & "00" & x"5a",
    "11" & x"3a" & "00" & x"ca",
    "10" & x"6a" & "10" & x"6a",
    "01" & x"6a" & "01" & x"6a",
    "11" & x"6a" & "00" & x"9a",
    "00" & x"ea" & "00" & x"ea",
    "10" & x"ea" & "01" & x"1a",
    "01" & x"ea" & "10" & x"1a",
    "10" & x"ba" & "01" & x"4a",
    "10" & x"76" & "01" & x"86",
    "01" & x"d6" & "10" & x"26",
    "10" & x"d6" & "01" & x"26",
    "11" & x"16" & "11" & x"16",
    "11" & x"56" & "00" & x"a6",
    "10" & x"96" & "10" & x"96",
    "01" & x"96" & "01" & x"96",
    "11" & x"86" & "00" & x"76",
    "11" & x"96" & "00" & x"66",
    "10" & x"56" & "10" & x"56",
    "01" & x"56" & "01" & x"56",
    "11" & x"46" & "11" & x"46",
    "00" & x"d6" & "00" & x"d6",
    "10" & x"c6" & "10" & x"c6",
    "01" & x"c6" & "01" & x"c6",
    "01" & x"76" & "10" & x"86",
    "01" & x"b6" & "10" & x"46",
    "10" & x"36" & "10" & x"36",
    "01" & x"36" & "01" & x"36",
    "11" & x"26" & "11" & x"26",
    "00" & x"b6" & "00" & x"b6",
    "10" & x"a6" & "10" & x"a6",
    "01" & x"a6" & "01" & x"a6",
    "11" & x"a6" & "00" & x"56",
    "11" & x"36" & "00" & x"c6",
    "10" & x"66" & "10" & x"66",
    "01" & x"66" & "01" & x"66",
    "11" & x"66" & "00" & x"96",
    "00" & x"e6" & "00" & x"e6",
    "10" & x"e6" & "01" & x"16",
    "01" & x"e6" & "10" & x"16",
    "10" & x"b6" & "01" & x"46",
    "10" & x"71" & "01" & x"8e",
    "01" & x"d1" & "10" & x"2e",
    "10" & x"d1" & "01" & x"2e",
    "11" & x"1e" & "11" & x"11",
    "11" & x"51" & "00" & x"ae",
    "10" & x"9e" & "10" & x"91",
    "01" & x"9e" & "01" & x"91",
    "11" & x"8e" & "00" & x"71",
    "11" & x"91" & "00" & x"6e",
    "10" & x"5e" & "10" & x"51",
    "01" & x"5e" & "01" & x"51",
    "11" & x"4e" & "11" & x"48",
    "00" & x"de" & "00" & x"d1",
    "10" & x"ce" & "10" & x"c8",
    "01" & x"ce" & "01" & x"c8",
    "01" & x"71" & "10" & x"8e",
    "01" & x"b1" & "10" & x"4e",
    "10" & x"37" & "10" & x"31",
    "01" & x"37" & "01" & x"31",
    "11" & x"2e" & "11" & x"21",
    "00" & x"b7" & "00" & x"b1",
    "10" & x"ae" & "10" & x"a1",
    "01" & x"ae" & "01" & x"a1",
    "11" & x"a1" & "00" & x"5e",
    "11" & x"31" & "00" & x"ce",
    "10" & x"6e" & "10" & x"61",
    "01" & x"6e" & "01" & x"61",
    "11" & x"61" & "00" & x"9e",
    "00" & x"ee" & "00" & x"e1",
    "10" & x"e1" & "01" & x"1e",
    "01" & x"e1" & "10" & x"1e",
    "10" & x"b1" & "01" & x"4e",
    "0011110100" & "1100001011",
    "0011111001" & "1100000110",
    "0011110101" & "1100001010",
    "0011110011" & "1100001100",
    "0011110010" & "1100001101",
    "0011111010" & "1100000101",
    "0011110110" & "1100001001",
    "0011111000" & "1100000111",
    "1110101000" & "0001010111",
    "1101101000" & "0010010111",
    "1011101000" & "0100010111",
    "0111101000" & "1000010111");

-- attribute ram_style : string;
-- attribute ram_style of ROM : signal is "block";


begin  -- behav


  clk_pra : process(clk) is
  begin
    if rising_edge(clk) then
      if rde_a = '1' then
        dout_a <= aRAM(to_integer(unsigned(address_a)));
      end if;
    end if;
  end process;

  clk_prb : process(clk) is
  begin
    if rising_edge(clk) then
      if rde_b = '1' then
        dout_b <= aRAM(to_integer(unsigned(address_b)));
      end if;
    end if;
  end process;
  

end behav;
